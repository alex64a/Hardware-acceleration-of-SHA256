`ifndef SHA256_SEQ_PKG_SV
 `define SHA256_SEQ_PKG_SV
package sha256_seq_pkg;
   import uvm_pkg::*;      // import the UVM library
 `include "uvm_macros.svh" // Include the UVM macros
  import sha256_agent_pkg::sha256_seq_item;
  import sha256_agent_pkg::sha256_sequencer;
 `include "sha256_base_seq.sv"
 `include "sha256_simple_seq.sv"
     endpackage 
`endif
